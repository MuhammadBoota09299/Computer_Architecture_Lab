module ALU (
    input logic [31:0]a,b,
    input logic [3:0]alu_op,
    output logic [31:0]result
);
    
endmodule