module napot (
    input logic [31:0] addr,addr_n,
    input logic [1:0]size,
    output logic napot_out
);
logic [4:0]position;
logic [31:0]ones,base,offset;

assign ones=~(32'b1 << position+1);
assign base=(addr_n & (ones));
assign offset=(32'h8<<position);
assign napot_out=(((base) + offset-1) >= (addr+size)) && (addr >= (base));



always_comb begin :priority_circuit
    casez (addr_n)  // casez allows ? for don't-care bits
        32'b???????????????????????????????0: position = 5'd0;
        32'b??????????????????????????????01: position = 5'd1;
        32'b?????????????????????????????011: position = 5'd2;
        32'b????????????????????????????0111: position = 5'd3;
        32'b???????????????????????????01111: position = 5'd4;
        32'b??????????????????????????011111: position = 5'd5;
        32'b?????????????????????????0111111: position = 5'd6;
        32'b????????????????????????01111111: position = 5'd7;
        32'b???????????????????????011111111: position = 5'd8;
        32'b??????????????????????0111111111: position = 5'd9;
        32'b?????????????????????01111111111: position = 5'd10;
        32'b????????????????????011111111111: position = 5'd11;
        32'b???????????????????0111111111111: position = 5'd12;
        32'b??????????????????01111111111111: position = 5'd13;
        32'b?????????????????011111111111111: position = 5'd14;
        32'b????????????????0111111111111111: position = 5'd15;
        32'b???????????????01111111111111111: position = 5'd16;
        32'b??????????????011111111111111111: position = 5'd17;
        32'b?????????????0111111111111111111: position = 5'd18;
        32'b????????????01111111111111111111: position = 5'd19;
        32'b???????????011111111111111111111: position = 5'd20;
        32'b??????????0111111111111111111111: position = 5'd21;
        32'b?????????01111111111111111111111: position = 5'd22;
        32'b????????011111111111111111111111: position = 5'd23;
        32'b???????0111111111111111111111111: position = 5'd24;
        32'b??????01111111111111111111111111: position = 5'd25;
        32'b?????011111111111111111111111111: position = 5'd26;
        32'b????0111111111111111111111111111: position = 5'd27;
        32'b???01111111111111111111111111111: position = 5'd28;
        32'b??011111111111111111111111111111: position = 5'd29;
        32'b?0111111111111111111111111111111: position = 5'd30;
        32'b01111111111111111111111111111111: position = 5'd31;
        default: position = 5'd0;  // When no bits are set
    endcase
end
    
endmodule