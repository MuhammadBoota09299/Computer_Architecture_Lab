module decoder (
    ports
);
    
endmodule