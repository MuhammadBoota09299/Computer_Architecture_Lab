module uart_tb ();
logic rx_bit,clock,reset;
log
endmodule