package single_cycle_processor
    typedef enum logic { 
        
     } opcodes;
endpackage